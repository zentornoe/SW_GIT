module cla_4bits (x,y,c_in,g_dot,p_dot,s); // 4bits Carry-Look-Ahead Adder

	input wire [3:0] x, y; // input operand : x, y
	input wire c_in; // input carry

	output wire g_dot, p_dot; // Group-generated carry, Group-propagated carry
	output wire [3:0] s; // output sum

	wire [3:0] g, p; // generated carry, propagated carry
	wire [3:0] c; // carry-look-ahead

	//coding here!!

    	/***********************
	//coding here!!
	//
	***********************/

endmodule
