module cla_16bits (x,y,c_in,s,c_out); // 16bits Carry-Look-Ahead Adder

	input wire [15:0] x, y; // input operand : x, y
	input wire c_in; // input carry

	output wire [15:0] s; // output sum
	output c_out; // output carry

	wire [3:0] g_dot, p_dot; // generated carry, propagated carry
	wire [3:0] c; // carry-look-ahead

	wire g_dot2, p_dot2; // Group-generated carry, Group-propagated carry

	//coding here!!

	/***********************
	//coding here!!
	//
	***********************/

	//coding here!!

endmodule

