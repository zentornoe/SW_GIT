module adder (x,y,c_in,g,p,s); // 1bit adder
	
	input wire x, y, c_in; // input operand : x, y  // input carry

	output wire g, p, s; // generated carry, propagated carry

	//coding here!!
	//coding here!!
	//coding here!!

endmodule
