module clag (g,p,c_in,c,g_dot,p_dot); // Carry-Look-Ahead Generator

	input wire [3:0] g, p; // generated carry, propagated carry
	input wire c_in; // input carry

	output wire [3:0] c; // carry-look-ahead
	output wire g_dot, p_dot; // generated carry, propagated carry

	/***********************
	//coding here!!
	//
	***********************/

	//coding here!!
	//coding here!!

endmodule

